library ieee;
use ieee.std_logic_1164.all;

package vector_pkg is
  type vector_t is array (natural range <>) of integer;
end package vector_pkg;
